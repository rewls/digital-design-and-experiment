`timescale 1 ns / 1 ns
`include "sha256.v"

`define test 512'h74657374800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020
`define SHA256 512'h53484132353680000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000030
`define META 512'h4d455441800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020
`define HDL 512'h48444c80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018

module top;

wire DONE;
wire [255:0] SHA256OUT;
reg CLK, nRST, START;
reg [511:0] SHA512IN;

sha256 test(DONE, SHA256OUT, CLK, nRST, START, SHA512IN);

initial begin
	CLK = 1'b0;
end

always begin
	#5 CLK = ~CLK;
end

initial begin
	nRST = 1'b0;
	#20 nRST = 1'b1;
end

initial begin
	START = 1'b0;
	#30 START = 1'b1;
	#10 START = 1'b0;
	#1010 $finish;
end

always @(START) begin
	if (START) begin
		SHA512IN = `test;
	end else begin
		SHA512IN = 512'h0;
	end
end

/*
initial
begin
    $dumpfile("test.vcd");
    $dumpvars(0, top);
end
*/

endmodule
